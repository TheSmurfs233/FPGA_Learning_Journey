module digit_rom_64x32(
    input [3:0] digit,      // 0-9数字编码
    input [7:0] row_addr,   // 行地址 0-63
    output reg [31:0] row_data // 32像素/行
);

// 每个数字64行x32列点阵数据
always @(*) begin
    case({digit, row_addr})
        // 数字0
        12'h000: row_data = 32'h00000000;
        12'h001: row_data = 32'h00000000;
        12'h002: row_data = 32'h00000000;
        12'h003: row_data = 32'h00000000;
        12'h004: row_data = 32'h00000000;
        12'h005: row_data = 32'h00000000;
        12'h006: row_data = 32'h00000000;
        12'h007: row_data = 32'h00000000;
        12'h008: row_data = 32'h00000000;
        12'h009: row_data = 32'h00000000;
        12'h00A: row_data = 32'h00000000;
        12'h00B: row_data = 32'h0007E000;
        12'h00C: row_data = 32'h001FF800;
        12'h00D: row_data = 32'h003C1E00;
        12'h00E: row_data = 32'h00700F00;
        12'h00F: row_data = 32'h00E00700;
        12'h010: row_data = 32'h01E00380;
        12'h011: row_data = 32'h03C003C0;
        12'h012: row_data = 32'h03C001C0;
        12'h013: row_data = 32'h078001E0;
        12'h014: row_data = 32'h078000E0;
        12'h015: row_data = 32'h070000E0;
        12'h016: row_data = 32'h0F0000F0;
        12'h017: row_data = 32'h0F0000F0;
        12'h018: row_data = 32'h0F0000F0;
        12'h019: row_data = 32'h0F000070;
        12'h01A: row_data = 32'h1E000078;
        12'h01B: row_data = 32'h1E000078;
        12'h01C: row_data = 32'h1E000078;
        12'h01D: row_data = 32'h1E000078;
        12'h01E: row_data = 32'h1E000078;
        12'h01F: row_data = 32'h1E000078;
        12'h020: row_data = 32'h1E000078;
        12'h021: row_data = 32'h1E000078;
        12'h022: row_data = 32'h1E000078;
        12'h023: row_data = 32'h1E000078;
        12'h024: row_data = 32'h1E000078;
        12'h025: row_data = 32'h1E000078;
        12'h026: row_data = 32'h1E000078;
        12'h027: row_data = 32'h1E000078;
        12'h028: row_data = 32'h0F000070;
        12'h029: row_data = 32'h0F0000F0;
        12'h02A: row_data = 32'h0F0000F0;
        12'h02B: row_data = 32'h0F0000F0;
        12'h02C: row_data = 32'h070000E0;
        12'h02D: row_data = 32'h078001E0;
        12'h02E: row_data = 32'h078001E0;
        12'h02F: row_data = 32'h03C001C0;
        12'h030: row_data = 32'h03C003C0;
        12'h031: row_data = 32'h01E00380;
        12'h032: row_data = 32'h00E00700;
        12'h033: row_data = 32'h00700F00;
        12'h034: row_data = 32'h003C1E00;
        12'h035: row_data = 32'h001FF800;
        12'h036: row_data = 32'h0007E000;
        12'h037: row_data = 32'h00000000;
        12'h038: row_data = 32'h00000000;
        12'h039: row_data = 32'h00000000;
        12'h03A: row_data = 32'h00000000;
        12'h03B: row_data = 32'h00000000;
        12'h03C: row_data = 32'h00000000;
        12'h03D: row_data = 32'h00000000;
        12'h03E: row_data = 32'h00000000;
        12'h03F: row_data = 32'h00000000;
        
        // 数字1
        12'h100: row_data = 32'h00000000;
        12'h101: row_data = 32'h00000000;
        12'h102: row_data = 32'h00000000;
        12'h103: row_data = 32'h00000000;
        12'h104: row_data = 32'h00000000;
        12'h105: row_data = 32'h00000000;
        12'h106: row_data = 32'h00000000;
        12'h107: row_data = 32'h00000000;
        12'h108: row_data = 32'h00000000;
        12'h109: row_data = 32'h00000000;
        12'h10A: row_data = 32'h00000000;
        12'h10B: row_data = 32'h00004000;
        12'h10C: row_data = 32'h0000C000;
        12'h10D: row_data = 32'h0001C000;
        12'h10E: row_data = 32'h0007C000;
        12'h10F: row_data = 32'h01FFC000;
        12'h110: row_data = 32'h01FFC000;
        12'h111: row_data = 32'h0007C000;
        12'h112: row_data = 32'h0003C000;
        12'h113: row_data = 32'h0003C000;
        12'h114: row_data = 32'h0003C000;
        12'h115: row_data = 32'h0003C000;
        12'h116: row_data = 32'h0003C000;
        12'h117: row_data = 32'h0003C000;
        12'h118: row_data = 32'h0003C000;
        12'h119: row_data = 32'h0003C000;
        12'h11A: row_data = 32'h0003C000;
        12'h11B: row_data = 32'h0003C000;
        12'h11C: row_data = 32'h0003C000;
        12'h11D: row_data = 32'h0003C000;
        12'h11E: row_data = 32'h0003C000;
        12'h11F: row_data = 32'h0003C000;
        12'h120: row_data = 32'h0003C000;
        12'h121: row_data = 32'h0003C000;
        12'h122: row_data = 32'h0003C000;
        12'h123: row_data = 32'h0003C000;
        12'h124: row_data = 32'h0003C000;
        12'h125: row_data = 32'h0003C000;
        12'h126: row_data = 32'h0003C000;
        12'h127: row_data = 32'h0003C000;
        12'h128: row_data = 32'h0003C000;
        12'h129: row_data = 32'h0003C000;
        12'h12A: row_data = 32'h0003C000;
        12'h12B: row_data = 32'h0003C000;
        12'h12C: row_data = 32'h0003C000;
        12'h12D: row_data = 32'h0003C000;
        12'h12E: row_data = 32'h0003C000;
        12'h12F: row_data = 32'h0003C000;
        12'h130: row_data = 32'h0003C000;
        12'h131: row_data = 32'h0003C000;
        12'h132: row_data = 32'h0003C000;
        12'h133: row_data = 32'h0007E000;
        12'h134: row_data = 32'h000FF000;
        12'h135: row_data = 32'h01FFFF80;
        12'h136: row_data = 32'h01FFFF80;
        12'h137: row_data = 32'h00000000;
        12'h138: row_data = 32'h00000000;
        12'h139: row_data = 32'h00000000;
        12'h13A: row_data = 32'h00000000;
        12'h13B: row_data = 32'h00000000;
        12'h13C: row_data = 32'h00000000;
        12'h13D: row_data = 32'h00000000;
        12'h13E: row_data = 32'h00000000;
        12'h13F: row_data = 32'h00000000;

        // 数字2
        12'h200: row_data = 32'h00000000;
        12'h201: row_data = 32'h00000000;
        12'h202: row_data = 32'h00000000;
        12'h203: row_data = 32'h00000000;
        12'h204: row_data = 32'h00000000;
        12'h205: row_data = 32'h00000000;
        12'h206: row_data = 32'h00000000;
        12'h207: row_data = 32'h00000000;
        12'h208: row_data = 32'h00000000;
        12'h209: row_data = 32'h00000000;
        12'h20A: row_data = 32'h00000000;
        12'h20B: row_data = 32'h000FF000;
        12'h20C: row_data = 32'h003FFE00;
        12'h20D: row_data = 32'h00F81F00;
        12'h20E: row_data = 32'h01E00780;
        12'h20F: row_data = 32'h03C003C0;
        12'h210: row_data = 32'h078001E0;
        12'h211: row_data = 32'h070001E0;
        12'h212: row_data = 32'h070000F0;
        12'h213: row_data = 32'h0F0000F0;
        12'h214: row_data = 32'h0F8000F0;
        12'h215: row_data = 32'h0F8000F0;
        12'h216: row_data = 32'h0FC000F0;
        12'h217: row_data = 32'h0FC000F0;
        12'h218: row_data = 32'h0FC000F0;
        12'h219: row_data = 32'h078001E0;
        12'h21A: row_data = 32'h000001E0;
        12'h21B: row_data = 32'h000001E0;
        12'h21C: row_data = 32'h000003C0;
        12'h21D: row_data = 32'h000003C0;
        12'h21E: row_data = 32'h00000780;
        12'h21F: row_data = 32'h00000F00;
        12'h220: row_data = 32'h00000E00;
        12'h221: row_data = 32'h00001C00;
        12'h222: row_data = 32'h00003800;
        12'h223: row_data = 32'h00007000;
        12'h224: row_data = 32'h0000E000;
        12'h225: row_data = 32'h0001C000;
        12'h226: row_data = 32'h00038000;
        12'h227: row_data = 32'h00070000;
        12'h228: row_data = 32'h000E0000;
        12'h229: row_data = 32'h001C0000;
        12'h22A: row_data = 32'h00380000;
        12'h22B: row_data = 32'h00700000;
        12'h22C: row_data = 32'h00E00030;
        12'h22D: row_data = 32'h01C00030;
        12'h22E: row_data = 32'h03800030;
        12'h22F: row_data = 32'h07800030;
        12'h230: row_data = 32'h07000060;
        12'h231: row_data = 32'h0E0000E0;
        12'h232: row_data = 32'h1C0001E0;
        12'h233: row_data = 32'h1FFFFFE0;
        12'h234: row_data = 32'h1FFFFFE0;
        12'h235: row_data = 32'h1FFFFFE0;
        12'h236: row_data = 32'h1FFFFFE0;
        12'h237: row_data = 32'h00000000;
        12'h238: row_data = 32'h00000000;
        12'h239: row_data = 32'h00000000;
        12'h23A: row_data = 32'h00000000;
        12'h23B: row_data = 32'h00000000;
        12'h23C: row_data = 32'h00000000;
        12'h23D: row_data = 32'h00000000;
        12'h23E: row_data = 32'h00000000;
        12'h23F: row_data = 32'h00000000;/*"2",0*/


        // 数字3
        12'h300: row_data = 32'h00000000;
        12'h301: row_data = 32'h00000000;
        12'h302: row_data = 32'h00000000;
        12'h303: row_data = 32'h00000000;
        12'h304: row_data = 32'h00000000;
        12'h305: row_data = 32'h00000000;
        12'h306: row_data = 32'h00000000;
        12'h307: row_data = 32'h00000000;
        12'h308: row_data = 32'h00000000;
        12'h309: row_data = 32'h00000000;
        12'h30A: row_data = 32'h00000000;
        12'h30B: row_data = 32'h000FE000;
        12'h30C: row_data = 32'h007FF800;
        12'h30D: row_data = 32'h00E07C00;
        12'h30E: row_data = 32'h01801E00;
        12'h30F: row_data = 32'h03000F00;
        12'h310: row_data = 32'h03000780;
        12'h311: row_data = 32'h07000780;
        12'h312: row_data = 32'h070007C0;
        12'h313: row_data = 32'h078003C0;
        12'h314: row_data = 32'h078003C0;
        12'h315: row_data = 32'h078003C0;
        12'h316: row_data = 32'h030003C0;
        12'h317: row_data = 32'h000003C0;
        12'h318: row_data = 32'h000003C0;
        12'h319: row_data = 32'h00000780;
        12'h31A: row_data = 32'h00000780;
        12'h31B: row_data = 32'h00000F00;
        12'h31C: row_data = 32'h00000E00;
        12'h31D: row_data = 32'h00003C00;
        12'h31E: row_data = 32'h0000F800;
        12'h31F: row_data = 32'h000FE000;
        12'h320: row_data = 32'h000FF800;
        12'h321: row_data = 32'h00007C00;
        12'h322: row_data = 32'h00000F00;
        12'h323: row_data = 32'h00000780;
        12'h324: row_data = 32'h000003C0;
        12'h325: row_data = 32'h000001C0;
        12'h326: row_data = 32'h000001E0;
        12'h327: row_data = 32'h000000E0;
        12'h328: row_data = 32'h000000F0;
        12'h329: row_data = 32'h000000F0;
        12'h32A: row_data = 32'h000000F0;
        12'h32B: row_data = 32'h038000F0;
        12'h32C: row_data = 32'h07C000F0;
        12'h32D: row_data = 32'h0FC000F0;
        12'h32E: row_data = 32'h0FC000F0;
        12'h32F: row_data = 32'h0FC001E0;
        12'h330: row_data = 32'h0F8001E0;
        12'h331: row_data = 32'h078003C0;
        12'h332: row_data = 32'h07800380;
        12'h333: row_data = 32'h03C00700;
        12'h334: row_data = 32'h01F01E00;
        12'h335: row_data = 32'h007FFC00;
        12'h336: row_data = 32'h001FE000;
        12'h337: row_data = 32'h00000000;
        12'h338: row_data = 32'h00000000;
        12'h339: row_data = 32'h00000000;
        12'h33A: row_data = 32'h00000000;
        12'h33B: row_data = 32'h00000000;
        12'h33C: row_data = 32'h00000000;
        12'h33D: row_data = 32'h00000000;
        12'h33E: row_data = 32'h00000000;
        12'h33F: row_data = 32'h00000000;/*"3",0*/


        // 数字4
        12'h400: row_data = 32'h00000000;
        12'h401: row_data = 32'h00000000;
        12'h402: row_data = 32'h00000000;
        12'h403: row_data = 32'h00000000;
        12'h404: row_data = 32'h00000000;
        12'h405: row_data = 32'h00000000;
        12'h406: row_data = 32'h00000000;
        12'h407: row_data = 32'h00000000;
        12'h408: row_data = 32'h00000000;
        12'h409: row_data = 32'h00000000;
        12'h40A: row_data = 32'h00000000;
        12'h40B: row_data = 32'h00000E00;
        12'h40C: row_data = 32'h00000E00;
        12'h40D: row_data = 32'h00001E00;
        12'h40E: row_data = 32'h00003E00;
        12'h40F: row_data = 32'h00003E00;
        12'h410: row_data = 32'h00007E00;
        12'h411: row_data = 32'h0000FE00;
        12'h412: row_data = 32'h0000DE00;
        12'h413: row_data = 32'h00019E00;
        12'h414: row_data = 32'h00039E00;
        12'h415: row_data = 32'h00031E00;
        12'h416: row_data = 32'h00071E00;
        12'h417: row_data = 32'h00061E00;
        12'h418: row_data = 32'h000C1E00;
        12'h419: row_data = 32'h001C1E00;
        12'h41A: row_data = 32'h00181E00;
        12'h41B: row_data = 32'h00301E00;
        12'h41C: row_data = 32'h00701E00;
        12'h41D: row_data = 32'h00601E00;
        12'h41E: row_data = 32'h00C01E00;
        12'h41F: row_data = 32'h01C01E00;
        12'h420: row_data = 32'h01801E00;
        12'h421: row_data = 32'h03001E00;
        12'h422: row_data = 32'h03001E00;
        12'h423: row_data = 32'h06001E00;
        12'h424: row_data = 32'h0E001E00;
        12'h425: row_data = 32'h0C001E00;
        12'h426: row_data = 32'h18001E00;
        12'h427: row_data = 32'h38001E00;
        12'h428: row_data = 32'h3FFFFFFC;
        12'h429: row_data = 32'h3FFFFFFC;
        12'h42A: row_data = 32'h00001E00;
        12'h42B: row_data = 32'h00001E00;
        12'h42C: row_data = 32'h00001E00;
        12'h42D: row_data = 32'h00001E00;
        12'h42E: row_data = 32'h00001E00;
        12'h42F: row_data = 32'h00001E00;
        12'h430: row_data = 32'h00001E00;
        12'h431: row_data = 32'h00001E00;
        12'h432: row_data = 32'h00001E00;
        12'h433: row_data = 32'h00001E00;
        12'h434: row_data = 32'h00003F00;
        12'h435: row_data = 32'h000FFFF8;
        12'h436: row_data = 32'h000FFFF8;
        12'h437: row_data = 32'h00000000;
        12'h438: row_data = 32'h00000000;
        12'h439: row_data = 32'h00000000;
        12'h43A: row_data = 32'h00000000;
        12'h43B: row_data = 32'h00000000;
        12'h43C: row_data = 32'h00000000;
        12'h43D: row_data = 32'h00000000;
        12'h43E: row_data = 32'h00000000;
        12'h43F: row_data = 32'h00000000;/*"4",0*/


        // 数字5
        12'h500: row_data = 32'h00000000;
        12'h501: row_data = 32'h00000000;
        12'h502: row_data = 32'h00000000;
        12'h503: row_data = 32'h00000000;
        12'h504: row_data = 32'h00000000;
        12'h505: row_data = 32'h00000000;
        12'h506: row_data = 32'h00000000;
        12'h507: row_data = 32'h00000000;
        12'h508: row_data = 32'h00000000;
        12'h509: row_data = 32'h00000000;
        12'h50A: row_data = 32'h00000000;
        12'h50B: row_data = 32'h01FFFFE0;
        12'h50C: row_data = 32'h01FFFFE0;
        12'h50D: row_data = 32'h01FFFFE0;
        12'h50E: row_data = 32'h01FFFFC0;
        12'h50F: row_data = 32'h01800000;
        12'h510: row_data = 32'h01800000;
        12'h511: row_data = 32'h01800000;
        12'h512: row_data = 32'h01800000;
        12'h513: row_data = 32'h01800000;
        12'h514: row_data = 32'h01800000;
        12'h515: row_data = 32'h01800000;
        12'h516: row_data = 32'h01800000;
        12'h517: row_data = 32'h01000000;
        12'h518: row_data = 32'h01000000;
        12'h519: row_data = 32'h03000000;
        12'h51A: row_data = 32'h0303F800;
        12'h51B: row_data = 32'h031FFE00;
        12'h51C: row_data = 32'h033FFF00;
        12'h51D: row_data = 32'h03781F80;
        12'h51E: row_data = 32'h036007C0;
        12'h51F: row_data = 32'h03C003C0;
        12'h520: row_data = 32'h038003E0;
        12'h521: row_data = 32'h038001E0;
        12'h522: row_data = 32'h000001E0;
        12'h523: row_data = 32'h000001F0;
        12'h524: row_data = 32'h000000F0;
        12'h525: row_data = 32'h000000F0;
        12'h526: row_data = 32'h000000F0;
        12'h527: row_data = 32'h000000F0;
        12'h528: row_data = 32'h000000F0;
        12'h529: row_data = 32'h000000F0;
        12'h52A: row_data = 32'h038000F0;
        12'h52B: row_data = 32'h07C000F0;
        12'h52C: row_data = 32'h0FC000F0;
        12'h52D: row_data = 32'h0FC000E0;
        12'h52E: row_data = 32'h0FC001E0;
        12'h52F: row_data = 32'h0F8001E0;
        12'h530: row_data = 32'h0F8001C0;
        12'h531: row_data = 32'h078003C0;
        12'h532: row_data = 32'h03800780;
        12'h533: row_data = 32'h01C00F00;
        12'h534: row_data = 32'h00F01E00;
        12'h535: row_data = 32'h007FFC00;
        12'h536: row_data = 32'h000FE000;
        12'h537: row_data = 32'h00000000;
        12'h538: row_data = 32'h00000000;
        12'h539: row_data = 32'h00000000;
        12'h53A: row_data = 32'h00000000;
        12'h53B: row_data = 32'h00000000;
        12'h53C: row_data = 32'h00000000;
        12'h53D: row_data = 32'h00000000;
        12'h53E: row_data = 32'h00000000;
        12'h53F: row_data = 32'h00000000;/*"5",0*/



        // 数字6
        12'h600: row_data = 32'h00000000;
        12'h601: row_data = 32'h00000000;
        12'h602: row_data = 32'h00000000;
        12'h603: row_data = 32'h00000000;
        12'h604: row_data = 32'h00000000;
        12'h605: row_data = 32'h00000000;
        12'h606: row_data = 32'h00000000;
        12'h607: row_data = 32'h00000000;
        12'h608: row_data = 32'h00000000;
        12'h609: row_data = 32'h00000000;
        12'h60A: row_data = 32'h00000000;
        12'h60B: row_data = 32'h0001FC00;
        12'h60C: row_data = 32'h0007FF00;
        12'h60D: row_data = 32'h001E0780;
        12'h60E: row_data = 32'h003803C0;
        12'h60F: row_data = 32'h007003E0;
        12'h610: row_data = 32'h00E003E0;
        12'h611: row_data = 32'h01C003E0;
        12'h612: row_data = 32'h038003E0;
        12'h613: row_data = 32'h038001C0;
        12'h614: row_data = 32'h07000000;
        12'h615: row_data = 32'h07000000;
        12'h616: row_data = 32'h07000000;
        12'h617: row_data = 32'h0F000000;
        12'h618: row_data = 32'h0F000000;
        12'h619: row_data = 32'h0E000000;
        12'h61A: row_data = 32'h0E000000;
        12'h61B: row_data = 32'h0E03F800;
        12'h61C: row_data = 32'h1E0FFF00;
        12'h61D: row_data = 32'h1E3FFF80;
        12'h61E: row_data = 32'h1E7C0FC0;
        12'h61F: row_data = 32'h1EF003E0;
        12'h620: row_data = 32'h1EE001E0;
        12'h621: row_data = 32'h1FC001F0;
        12'h622: row_data = 32'h1F8000F0;
        12'h623: row_data = 32'h1F0000F0;
        12'h624: row_data = 32'h1F000078;
        12'h625: row_data = 32'h1E000078;
        12'h626: row_data = 32'h1E000078;
        12'h627: row_data = 32'h1E000078;
        12'h628: row_data = 32'h1E000078;
        12'h629: row_data = 32'h1E000078;
        12'h62A: row_data = 32'h0E000078;
        12'h62B: row_data = 32'h0F000078;
        12'h62C: row_data = 32'h0F000078;
        12'h62D: row_data = 32'h0F000070;
        12'h62E: row_data = 32'h070000F0;
        12'h62F: row_data = 32'h078000F0;
        12'h630: row_data = 32'h03C000E0;
        12'h631: row_data = 32'h03C001E0;
        12'h632: row_data = 32'h01E001C0;
        12'h633: row_data = 32'h00F00380;
        12'h634: row_data = 32'h007C0F00;
        12'h635: row_data = 32'h003FFE00;
        12'h636: row_data = 32'h0007F000;
        12'h637: row_data = 32'h00000000;
        12'h638: row_data = 32'h00000000;
        12'h639: row_data = 32'h00000000;
        12'h63A: row_data = 32'h00000000;
        12'h63B: row_data = 32'h00000000;
        12'h63C: row_data = 32'h00000000;
        12'h63D: row_data = 32'h00000000;
        12'h63E: row_data = 32'h00000000;
        12'h63F: row_data = 32'h00000000;/*"6",0*/



        // 数字7
        12'h700: row_data = 32'h00000000;
        12'h701: row_data = 32'h00000000;
        12'h702: row_data = 32'h00000000;
        12'h703: row_data = 32'h00000000;
        12'h704: row_data = 32'h00000000;
        12'h705: row_data = 32'h00000000;
        12'h706: row_data = 32'h00000000;
        12'h707: row_data = 32'h00000000;
        12'h708: row_data = 32'h00000000;
        12'h709: row_data = 32'h00000000;
        12'h70A: row_data = 32'h00000000;
        12'h70B: row_data = 32'h03FFFFF0;
        12'h70C: row_data = 32'h07FFFFF0;
        12'h70D: row_data = 32'h07FFFFF0;
        12'h70E: row_data = 32'h07FFFFE0;
        12'h70F: row_data = 32'h07C000C0;
        12'h710: row_data = 32'h070000C0;
        12'h711: row_data = 32'h06000180;
        12'h712: row_data = 32'h06000180;
        12'h713: row_data = 32'h0C000300;
        12'h714: row_data = 32'h0C000300;
        12'h715: row_data = 32'h0C000600;
        12'h716: row_data = 32'h00000600;
        12'h717: row_data = 32'h00000C00;
        12'h718: row_data = 32'h00001C00;
        12'h719: row_data = 32'h00001800;
        12'h71A: row_data = 32'h00003800;
        12'h71B: row_data = 32'h00003800;
        12'h71C: row_data = 32'h00003000;
        12'h71D: row_data = 32'h00007000;
        12'h71E: row_data = 32'h00007000;
        12'h71F: row_data = 32'h0000E000;
        12'h720: row_data = 32'h0000E000;
        12'h721: row_data = 32'h0001E000;
        12'h722: row_data = 32'h0001C000;
        12'h723: row_data = 32'h0003C000;
        12'h724: row_data = 32'h0003C000;
        12'h725: row_data = 32'h00038000;
        12'h726: row_data = 32'h00078000;
        12'h727: row_data = 32'h00078000;
        12'h728: row_data = 32'h00078000;
        12'h729: row_data = 32'h000F8000;
        12'h72A: row_data = 32'h000F8000;
        12'h72B: row_data = 32'h000F8000;
        12'h72C: row_data = 32'h000F8000;
        12'h72D: row_data = 32'h000F8000;
        12'h72E: row_data = 32'h001F8000;
        12'h72F: row_data = 32'h001F8000;
        12'h730: row_data = 32'h001F8000;
        12'h731: row_data = 32'h001F8000;
        12'h732: row_data = 32'h001F8000;
        12'h733: row_data = 32'h001F8000;
        12'h734: row_data = 32'h001F8000;
        12'h735: row_data = 32'h001F8000;
        12'h736: row_data = 32'h000F0000;
        12'h737: row_data = 32'h00000000;
        12'h738: row_data = 32'h00000000;
        12'h739: row_data = 32'h00000000;
        12'h73A: row_data = 32'h00000000;
        12'h73B: row_data = 32'h00000000;
        12'h73C: row_data = 32'h00000000;
        12'h73D: row_data = 32'h00000000;
        12'h73E: row_data = 32'h00000000;
        12'h73F: row_data = 32'h00000000;/*"7",0*/


        // 数字8
        12'h800: row_data = 32'h00000000;
        12'h801: row_data = 32'h00000000;
        12'h802: row_data = 32'h00000000;
        12'h803: row_data = 32'h00000000;
        12'h804: row_data = 32'h00000000;
        12'h805: row_data = 32'h00000000;
        12'h806: row_data = 32'h00000000;
        12'h807: row_data = 32'h00000000;
        12'h808: row_data = 32'h00000000;
        12'h809: row_data = 32'h00000000;
        12'h80A: row_data = 32'h00000000;
        12'h80B: row_data = 32'h000FF000;
        12'h80C: row_data = 32'h007FFE00;
        12'h80D: row_data = 32'h00F81F00;
        12'h80E: row_data = 32'h01E00780;
        12'h80F: row_data = 32'h03C003C0;
        12'h810: row_data = 32'h078001E0;
        12'h811: row_data = 32'h078001E0;
        12'h812: row_data = 32'h0F0000F0;
        12'h813: row_data = 32'h0F0000F0;
        12'h814: row_data = 32'h0F0000F0;
        12'h815: row_data = 32'h0F0000F0;
        12'h816: row_data = 32'h0F0000F0;
        12'h817: row_data = 32'h0F8000F0;
        12'h818: row_data = 32'h0F8000E0;
        12'h819: row_data = 32'h07C001E0;
        12'h81A: row_data = 32'h07E001C0;
        12'h81B: row_data = 32'h03F003C0;
        12'h81C: row_data = 32'h01FC0780;
        12'h81D: row_data = 32'h00FF0E00;
        12'h81E: row_data = 32'h007FDC00;
        12'h81F: row_data = 32'h001FF000;
        12'h820: row_data = 32'h003FF800;
        12'h821: row_data = 32'h00F1FE00;
        12'h822: row_data = 32'h01E07F00;
        12'h823: row_data = 32'h03C03F80;
        12'h824: row_data = 32'h07801FC0;
        12'h825: row_data = 32'h078007C0;
        12'h826: row_data = 32'h0F0003E0;
        12'h827: row_data = 32'h0F0003E0;
        12'h828: row_data = 32'h1E0001F0;
        12'h829: row_data = 32'h1E0001F0;
        12'h82A: row_data = 32'h1E0000F0;
        12'h82B: row_data = 32'h1E0000F0;
        12'h82C: row_data = 32'h1E0000F0;
        12'h82D: row_data = 32'h1E0000F0;
        12'h82E: row_data = 32'h1E0000F0;
        12'h82F: row_data = 32'h0F0000E0;
        12'h830: row_data = 32'h0F0001E0;
        12'h831: row_data = 32'h078001C0;
        12'h832: row_data = 32'h078003C0;
        12'h833: row_data = 32'h03E00780;
        12'h834: row_data = 32'h00F81F00;
        12'h835: row_data = 32'h007FFC00;
        12'h836: row_data = 32'h000FF000;
        12'h837: row_data = 32'h00000000;
        12'h838: row_data = 32'h00000000;
        12'h839: row_data = 32'h00000000;
        12'h83A: row_data = 32'h00000000;
        12'h83B: row_data = 32'h00000000;
        12'h83C: row_data = 32'h00000000;
        12'h83D: row_data = 32'h00000000;
        12'h83E: row_data = 32'h00000000;
        12'h83F: row_data = 32'h00000000;

        
        // 数字9
        12'h900: row_data = 32'h00000000;
        12'h901: row_data = 32'h00000000;
        12'h902: row_data = 32'h00000000;
        12'h903: row_data = 32'h00000000;
        12'h904: row_data = 32'h00000000;
        12'h905: row_data = 32'h00000000;
        12'h906: row_data = 32'h00000000;
        12'h907: row_data = 32'h00000000;
        12'h908: row_data = 32'h00000000;
        12'h909: row_data = 32'h00000000;
        12'h90A: row_data = 32'h00000000;
        12'h90B: row_data = 32'h001FE000;
        12'h90C: row_data = 32'h007FF800;
        12'h90D: row_data = 32'h00F03C00;
        12'h90E: row_data = 32'h01E00E00;
        12'h90F: row_data = 32'h03C00700;
        12'h910: row_data = 32'h07800380;
        12'h911: row_data = 32'h07000380;
        12'h912: row_data = 32'h0F0001C0;
        12'h913: row_data = 32'h0F0001C0;
        12'h914: row_data = 32'h0E0001E0;
        12'h915: row_data = 32'h1E0000E0;
        12'h916: row_data = 32'h1E0000E0;
        12'h917: row_data = 32'h1E0000E0;
        12'h918: row_data = 32'h1E0000F0;
        12'h919: row_data = 32'h1E0000F0;
        12'h91A: row_data = 32'h1E0000F0;
        12'h91B: row_data = 32'h1E0000F0;
        12'h91C: row_data = 32'h1E0000F0;
        12'h91D: row_data = 32'h1E0001F0;
        12'h91E: row_data = 32'h1F0001F0;
        12'h91F: row_data = 32'h0F0003F0;
        12'h920: row_data = 32'h0F8006F0;
        12'h921: row_data = 32'h0F800EF0;
        12'h922: row_data = 32'h07C01CF0;
        12'h923: row_data = 32'h03F07CF0;
        12'h924: row_data = 32'h01FFF8F0;
        12'h925: row_data = 32'h00FFE0F0;
        12'h926: row_data = 32'h003F81E0;
        12'h927: row_data = 32'h000001E0;
        12'h928: row_data = 32'h000001E0;
        12'h929: row_data = 32'h000001E0;
        12'h92A: row_data = 32'h000001C0;
        12'h92B: row_data = 32'h000003C0;
        12'h92C: row_data = 32'h000003C0;
        12'h92D: row_data = 32'h00000380;
        12'h92E: row_data = 32'h03800780;
        12'h92F: row_data = 32'h07C00700;
        12'h930: row_data = 32'h07C00F00;
        12'h931: row_data = 32'h07C00E00;
        12'h932: row_data = 32'h07C01C00;
        12'h933: row_data = 32'h03C03800;
        12'h934: row_data = 32'h03E0F000;
        12'h935: row_data = 32'h01FFE000;
        12'h936: row_data = 32'h003F0000;
        12'h937: row_data = 32'h00000000;
        12'h938: row_data = 32'h00000000;
        12'h939: row_data = 32'h00000000;
        12'h93A: row_data = 32'h00000000;
        12'h93B: row_data = 32'h00000000;
        12'h93C: row_data = 32'h00000000;
        12'h93D: row_data = 32'h00000000;
        12'h93E: row_data = 32'h00000000;
        12'h93F: row_data = 32'h00000000;

        default: row_data = 32'h0000;
    endcase
end

endmodule