module vga_image_gen (
    input  vga_clk,
    input  rst_n,
    input [9:0] pix_x,
    input [9:0] pix_y,  
    output reg [15:0] pix_data
);

//parameter definition
parameter CHAR_B_H= 10'd63 ; //字符开始X轴坐标
parameter CHAR_B_V= 10'd208 ; //字符开始Y轴坐标
parameter CHAR_W = 10'd512 ; //字符宽度
parameter CHAR_H = 10'd64 ; //字符高度
parameter BLACK = 16'h0000; //黑色
parameter WHITE = 16'hFFFF; //白色
parameter GOLDEN = 16'hFEC0; //金色

//wire definition
wire [9:0] char_x;   //字符X轴坐标
wire [9:0] char_y;   //字符Y轴坐标

//reg define
reg [0:511] char [63:0] ; //字符数据


/****** main logic ******/

//字符显示坐标
assign char_x = ((pix_x >= CHAR_B_H) && (pix_y>= CHAR_B_V) && (pix_x <= (CHAR_B_H + CHAR_W)) && (pix_y <= (CHAR_B_V + CHAR_H) )) ? (pix_x - CHAR_B_H - 1'b1):10'h3FF;
assign char_y = ((pix_x >= CHAR_B_H) && (pix_y>= CHAR_B_V) && (pix_x <= (CHAR_B_H + CHAR_W)) && (pix_y <= (CHAR_B_V + CHAR_H) )) ? (pix_y - CHAR_B_V - 1'b1):10'h3FF;

//pix_data:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
always @(posedge vga_clk ,negedge rst_n) begin
    if (rst_n == 1'b0) begin
        pix_data <= 16'h0000;
    end 
    else begin
        if ((char_x == 10'h3FF) || (char_y == 10'h3FF)) begin
            pix_data <= BLACK;
        end 
        else begin
            pix_data <= char[char_y][char_x] ? GOLDEN : BLACK;
        end
    end
end

//char:字符数据初始化
always @(posedge vga_clk ) begin
    char[0]  <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[1]  <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[2]  <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[3]  <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[4]  <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[5]  <= 512'h0000001E000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000180000000000000000000000;
    char[6]  <= 512'h0000001F8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001F000000000000003C000000;
    char[7]  <= 512'h0000001FE0000000000000000000000000000000000000000000000E000000000000000003E000000000000018000000000000001F800000000000003F000000;
    char[8]  <= 512'h0000000FE00000000000000000000000000000000000000000000007E000000000000001FFF800000000F0001E000000000000000F800000000000001E000000;
    char[9]  <= 512'h0000000FE00000000000000000000000000000000000000000000003E0000000000003FFC3F000000000FC001F000000000000000F800000000000003C000000;
    char[10] <= 512'h0000001FC000000000003E00000E0000000000000000000000000003E0000000000001F003C0000000007C001E000000000000000F800000000000003C380000;
    char[11] <= 512'h0000001F800000000000FF8001FF8000000000000E00000000000003C000C0000000000007800000000078003C000000000003C0070000000000000038FF0000;
    char[12] <= 512'h0000001F0000000000F7FF00FF07E000000000007F80000000070003C001F000000000781E000000000078003F000000000001F007000000000000007FFF0000;
    char[13] <= 512'h0000003E003C0000007F1EFF7807F0000000001FFFE000000007E003C001F8000000000FFC0000000000780079800000000001F80700000000007C00E03E0000;
    char[14] <= 512'h0000003E07FFC000003C3C703C07E0000001FFFFFFF000000003F003C003F00000000001FC0000000000700070E00000000000F00700F00000C7FF01C0780000;
    char[15] <= 512'h0000007DFFFFE000003C38703C07C0000000FFF81FE000000001F003C007800000000003FF00000000007000F0700000000000F00707F80000FFFF0180F00000;
    char[16] <= 512'h00000FFFFFFFC000003C30303C07800000001C001F8000000000F0038C0E00000000000F8F80000000007000E03C0000000000F007FFF80000783E0300E00000;
    char[17] <= 512'h001FFFFFFFC00000003C70303FE78000000000001E00000000000003FDF800000000003E01C0000000007001C01E0000000000F007FE000000781C0601800000;
    char[18] <= 512'h000FFFFC00000000001C6033FF870000000000003C0000000000001FF1E00000000001F0001F8000000070038007800000000FF00700000000781C0803000000;
    char[19] <= 512'h0001C1E000000000001C6011F80F0000000000003C000000000001FFC0E000000000000003FFC000000070070003E0000003FFF00700000000781C00060F8000;
    char[20] <= 512'h000003E000000000001C6018380E00000007800038000000000001FF80E000000000003C1F8F000000006F0F0001F800001FF8700700000000381C000DFFE000;
    char[21] <= 512'h000007CFC0000000001C3018380E00000003C000780000000000000380E01F0000003FFF001E00000001FF8E03E0FE00000780700700000000381C007F03F000;
    char[22] <= 512'h00000F87E0000000001C3018781E00000003E000780000000000000380E1FF8000007F1F201C0000003FFE183FE07FE0000000700700000000381C7FCC03F000;
    char[23] <= 512'h00000F07E0000000001C18187FFC00000003E000FC0000000003C0039CFFFC000000001C3E38000001FFE031FF003FFC000000700703F00000381C780E03C000;
    char[24] <= 512'h00001F03E0000000001C1C0FFFFC00000003E03FFC000000000FF003F8FF80000000303807F000000001E06000000FF000000070077FF00000381C380E038000;
    char[25] <= 512'h00003E03E0000000001DFC0FF81800000001FFFF8000000000FFF003E0E1C00000001C7001FC00000001E180000600000000007007FF8000003BDC1C0C070000;
    char[26] <= 512'h00007C03E0000000001CFC0C380000000001FF80000000000071E00780E1C000000007E007BF00000003E3000007800000000FF007000000003FDC1C0C060000;
    char[27] <= 512'h0000F803E7FE0000001C3C00380000000001C000000000000001C03F80C1C000000003C01E0FC000000760000003C0000003FFF00700000000381C1C0C3F0000;
    char[28] <= 512'h0003F007FFFF0000001C1C003801F0000001C00000000000000380FB80C1C000000007F07803C00000066001C103C0000003F8700700000000381C0C1FFF0000;
    char[29] <= 512'h000FFFFFFF800000001C0C00387FFE000001800000000000000383F381C1C00000001E780000C000000EFC7FE1838000000000700700000000381C0FFF000000;
    char[30] <= 512'h000FFFE3E0000000001C00003FF03F00000380000000000000030FC381C1C00000003839C0000000001CFE30E1C18000000000700700000000381C0FB8000000;
    char[31] <= 512'h0007E003E0000000001C060FFC003E00000380000000000000030F8381C1C0000000C001E000FF800018EE30E1C18000000000700700000000381C0438000000;
    char[32] <= 512'h00078003E0000000001C07F838003E000003800000000200000382038381C00000000000E1FFFFC00038E030E1C18000000000700700FE0000381C0073800000;
    char[33] <= 512'h00000003E0000000001C038038003C000003800000000200000380038381C00000000003FFFFFFC00070E030E1C18000000007F0070FFF8000381C0073C00000;
    char[34] <= 512'h00003003E0000000003C038038703C0000038000000002000001C0078301C00000001FFFE000000000E0E03FE1C1C0000001FFF007FFFF8000381C00E3C00000;
    char[35] <= 512'h00007003E0FC0000003C038038383C0000038000000006000001C0078601C000007FFF8FF800000001C0E030E1C1C000007FFC7007FFC00000781C01C3800000;
    char[36] <= 512'h0000F003E07F8000003C038039FC3C0000038000000006000000C03F8E01C000003FC00EFC0000000300E030E1C1C000007FC07007000000007BFC03C3800010;
    char[37] <= 512'h0001F003E03FE000003C0380FE1C3C000003800000000F000000C01F0C01C0000000001CEF0000000600E070E1C1C000000000F007000000007FDC0783800010;
    char[38] <= 512'h0003F003E01FF000003C039FE01C3C000003C00000000F000000C00F1801C0000000003CE38000000800E07FE1C1C000000000F00700000000381C0F03800018;
    char[39] <= 512'h0007F003E00FF800003C038F00003C000001E00000001F00001FF8060001C00000000078E1E000000001E060E181C000000000F0070000000038181E03800018;
    char[40] <= 512'h000FE003E007FC00007C038000003C000001F00000007F0001FFFF8000018000000001E0E0F800000001C060E001C000000000F00F0000000000003C03800038;
    char[41] <= 512'h001FC003E003FC00007C0380000078000000FC000003FF0001F807FC00018000000003C0E07E00000001C0E0E001C000000001F00F0000000000007003800038;
    char[42] <= 512'h001F8003E001FC00007803800000780000007FC0007FFF000060007FE001800000000780E03FC0000001C0E0E001C000000001F00F000000000001E00380007C;
    char[43] <= 512'h001F0003E000FC0000780380001FF80000001FFFFFFFFC0000000007FFC0000000001E00E00FFC000003C0C0E001C000000001E00F0000000000078001C000FC;
    char[44] <= 512'h001E01FFE000380000780380000FF000000003FFFFFFC00000000000FFFFFFFC00007C00E007FFE00003C0C0E003C000000001E00F00000000000E0001F007FC;
    char[45] <= 512'h001800FFE0000000007801800007F0000000001FFFF00000000000000FFFFFF00001E001E001FFF80001C00FE023C000000000E00F0000000000100000FFFFF8;
    char[46] <= 512'h0000007FE0000000003000000003E00000000000000000000000000001FFFE0000078001E0007E000001C007C03FC000000000000F00000000000000007FFFE0;
    char[47] <= 512'h0000003FC0000000000000000003C000000000000000000000000000001FE000001C0001E000000000008003C00F8000000000000F00000000000000000FFE00;
    char[48] <= 512'h0000000F8000000000000000000100000000000000000000000000000000000000000000E00000000000000180078000000000000F0000000000000000000000;
    char[49] <= 512'h000000070000000000000000000000000000000000000000000000000000000000000000E0000000000000000007000000000000060000000000000000000000;
    char[50] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000040000000000000000002000000000000000000000000000000000000;
    char[51] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[52] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[53] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[54] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[55] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[56] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[57] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[58] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[59] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[60] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[61] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[62] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    char[63] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end
endmodule